// Gshare Predictor

module gshare();

endmodule