// Branch Prediction Unit

module BPU(in_PC, in_hit, out_predict);

endmodule