// Bimodal Predictor

module bimodal();

endmodule