// Branch Prediction Unit

module BPU(in_PC, in_hit, out_predict);
    input   in_PC, in_hit;
    output  out_predict;
endmodule