// Square-root Normaliser
module Sqrt_Norm(in_Exp, in_Mant, out_Exp, out_Mant);
    input   [7:0]   in_Exp;
    input   [253:0] in_Mant;

    output reg [7:0]   out_Exp;
    output reg [253:0]  out_Mant;

    always @ (*) begin
        if (in_Mant[253]) begin out_Exp = in_Exp + 8'd126; out_Mant = in_Mant >> 126; end
        else if (in_Mant[252]) begin out_Exp = in_Exp + 8'd125; out_Mant = in_Mant >> 125; end
        else if (in_Mant[251]) begin out_Exp = in_Exp + 8'd124; out_Mant = in_Mant >> 124; end
        else if (in_Mant[250]) begin out_Exp = in_Exp + 8'd123; out_Mant = in_Mant >> 123; end
        else if (in_Mant[249]) begin out_Exp = in_Exp + 8'd122; out_Mant = in_Mant >> 122; end
        else if (in_Mant[248]) begin out_Exp = in_Exp + 8'd121; out_Mant = in_Mant >> 121; end
        else if (in_Mant[247]) begin out_Exp = in_Exp + 8'd120; out_Mant = in_Mant >> 120; end
        else if (in_Mant[246]) begin out_Exp = in_Exp + 8'd119; out_Mant = in_Mant >> 119; end
        else if (in_Mant[245]) begin out_Exp = in_Exp + 8'd118; out_Mant = in_Mant >> 118; end
        else if (in_Mant[244]) begin out_Exp = in_Exp + 8'd117; out_Mant = in_Mant >> 117; end
        else if (in_Mant[243]) begin out_Exp = in_Exp + 8'd116; out_Mant = in_Mant >> 116; end
        else if (in_Mant[242]) begin out_Exp = in_Exp + 8'd115; out_Mant = in_Mant >> 115; end
        else if (in_Mant[241]) begin out_Exp = in_Exp + 8'd114; out_Mant = in_Mant >> 114; end
        else if (in_Mant[240]) begin out_Exp = in_Exp + 8'd113; out_Mant = in_Mant >> 113; end
        else if (in_Mant[239]) begin out_Exp = in_Exp + 8'd112; out_Mant = in_Mant >> 112; end
        else if (in_Mant[238]) begin out_Exp = in_Exp + 8'd111; out_Mant = in_Mant >> 111; end
        else if (in_Mant[237]) begin out_Exp = in_Exp + 8'd110; out_Mant = in_Mant >> 110; end
        else if (in_Mant[236]) begin out_Exp = in_Exp + 8'd109; out_Mant = in_Mant >> 109; end
        else if (in_Mant[235]) begin out_Exp = in_Exp + 8'd108; out_Mant = in_Mant >> 108; end
        else if (in_Mant[234]) begin out_Exp = in_Exp + 8'd107; out_Mant = in_Mant >> 107; end
        else if (in_Mant[233]) begin out_Exp = in_Exp + 8'd106; out_Mant = in_Mant >> 106; end
        else if (in_Mant[232]) begin out_Exp = in_Exp + 8'd105; out_Mant = in_Mant >> 105; end
        else if (in_Mant[231]) begin out_Exp = in_Exp + 8'd104; out_Mant = in_Mant >> 104; end
        else if (in_Mant[230]) begin out_Exp = in_Exp + 8'd103; out_Mant = in_Mant >> 103; end
        else if (in_Mant[229]) begin out_Exp = in_Exp + 8'd102; out_Mant = in_Mant >> 102; end
        else if (in_Mant[228]) begin out_Exp = in_Exp + 8'd101; out_Mant = in_Mant >> 101; end
        else if (in_Mant[227]) begin out_Exp = in_Exp + 8'd100; out_Mant = in_Mant >> 100; end
        else if (in_Mant[226]) begin out_Exp = in_Exp + 8'd99; out_Mant = in_Mant >> 99; end
        else if (in_Mant[225]) begin out_Exp = in_Exp + 8'd98; out_Mant = in_Mant >> 98; end
        else if (in_Mant[224]) begin out_Exp = in_Exp + 8'd97; out_Mant = in_Mant >> 97; end
        else if (in_Mant[223]) begin out_Exp = in_Exp + 8'd96; out_Mant = in_Mant >> 96; end
        else if (in_Mant[222]) begin out_Exp = in_Exp + 8'd95; out_Mant = in_Mant >> 95; end
        else if (in_Mant[221]) begin out_Exp = in_Exp + 8'd94; out_Mant = in_Mant >> 94; end
        else if (in_Mant[220]) begin out_Exp = in_Exp + 8'd93; out_Mant = in_Mant >> 93; end
        else if (in_Mant[219]) begin out_Exp = in_Exp + 8'd92; out_Mant = in_Mant >> 92; end
        else if (in_Mant[218]) begin out_Exp = in_Exp + 8'd91; out_Mant = in_Mant >> 91; end
        else if (in_Mant[217]) begin out_Exp = in_Exp + 8'd90; out_Mant = in_Mant >> 90; end
        else if (in_Mant[216]) begin out_Exp = in_Exp + 8'd89; out_Mant = in_Mant >> 89; end
        else if (in_Mant[215]) begin out_Exp = in_Exp + 8'd88; out_Mant = in_Mant >> 88; end
        else if (in_Mant[214]) begin out_Exp = in_Exp + 8'd87; out_Mant = in_Mant >> 87; end
        else if (in_Mant[213]) begin out_Exp = in_Exp + 8'd86; out_Mant = in_Mant >> 86; end
        else if (in_Mant[212]) begin out_Exp = in_Exp + 8'd85; out_Mant = in_Mant >> 85; end
        else if (in_Mant[211]) begin out_Exp = in_Exp + 8'd84; out_Mant = in_Mant >> 84; end
        else if (in_Mant[210]) begin out_Exp = in_Exp + 8'd83; out_Mant = in_Mant >> 83; end
        else if (in_Mant[209]) begin out_Exp = in_Exp + 8'd82; out_Mant = in_Mant >> 82; end
        else if (in_Mant[208]) begin out_Exp = in_Exp + 8'd81; out_Mant = in_Mant >> 81; end
        else if (in_Mant[207]) begin out_Exp = in_Exp + 8'd80; out_Mant = in_Mant >> 80; end
        else if (in_Mant[206]) begin out_Exp = in_Exp + 8'd79; out_Mant = in_Mant >> 79; end
        else if (in_Mant[205]) begin out_Exp = in_Exp + 8'd78; out_Mant = in_Mant >> 78; end
        else if (in_Mant[204]) begin out_Exp = in_Exp + 8'd77; out_Mant = in_Mant >> 77; end
        else if (in_Mant[203]) begin out_Exp = in_Exp + 8'd76; out_Mant = in_Mant >> 76; end
        else if (in_Mant[202]) begin out_Exp = in_Exp + 8'd75; out_Mant = in_Mant >> 75; end
        else if (in_Mant[201]) begin out_Exp = in_Exp + 8'd74; out_Mant = in_Mant >> 74; end
        else if (in_Mant[200]) begin out_Exp = in_Exp + 8'd73; out_Mant = in_Mant >> 73; end
        else if (in_Mant[199]) begin out_Exp = in_Exp + 8'd72; out_Mant = in_Mant >> 72; end
        else if (in_Mant[198]) begin out_Exp = in_Exp + 8'd71; out_Mant = in_Mant >> 71; end
        else if (in_Mant[197]) begin out_Exp = in_Exp + 8'd70; out_Mant = in_Mant >> 70; end
        else if (in_Mant[196]) begin out_Exp = in_Exp + 8'd69; out_Mant = in_Mant >> 69; end
        else if (in_Mant[195]) begin out_Exp = in_Exp + 8'd68; out_Mant = in_Mant >> 68; end
        else if (in_Mant[194]) begin out_Exp = in_Exp + 8'd67; out_Mant = in_Mant >> 67; end
        else if (in_Mant[193]) begin out_Exp = in_Exp + 8'd66; out_Mant = in_Mant >> 66; end
        else if (in_Mant[192]) begin out_Exp = in_Exp + 8'd65; out_Mant = in_Mant >> 65; end
        else if (in_Mant[191]) begin out_Exp = in_Exp + 8'd64; out_Mant = in_Mant >> 64; end
        else if (in_Mant[190]) begin out_Exp = in_Exp + 8'd63; out_Mant = in_Mant >> 63; end
        else if (in_Mant[189]) begin out_Exp = in_Exp + 8'd62; out_Mant = in_Mant >> 62; end
        else if (in_Mant[188]) begin out_Exp = in_Exp + 8'd61; out_Mant = in_Mant >> 61; end
        else if (in_Mant[187]) begin out_Exp = in_Exp + 8'd60; out_Mant = in_Mant >> 60; end
        else if (in_Mant[186]) begin out_Exp = in_Exp + 8'd59; out_Mant = in_Mant >> 59; end
        else if (in_Mant[185]) begin out_Exp = in_Exp + 8'd58; out_Mant = in_Mant >> 58; end
        else if (in_Mant[184]) begin out_Exp = in_Exp + 8'd57; out_Mant = in_Mant >> 57; end
        else if (in_Mant[183]) begin out_Exp = in_Exp + 8'd56; out_Mant = in_Mant >> 56; end
        else if (in_Mant[182]) begin out_Exp = in_Exp + 8'd55; out_Mant = in_Mant >> 55; end
        else if (in_Mant[181]) begin out_Exp = in_Exp + 8'd54; out_Mant = in_Mant >> 54; end
        else if (in_Mant[180]) begin out_Exp = in_Exp + 8'd53; out_Mant = in_Mant >> 53; end
        else if (in_Mant[179]) begin out_Exp = in_Exp + 8'd52; out_Mant = in_Mant >> 52; end
        else if (in_Mant[178]) begin out_Exp = in_Exp + 8'd51; out_Mant = in_Mant >> 51; end
        else if (in_Mant[177]) begin out_Exp = in_Exp + 8'd50; out_Mant = in_Mant >> 50; end
        else if (in_Mant[176]) begin out_Exp = in_Exp + 8'd49; out_Mant = in_Mant >> 49; end
        else if (in_Mant[175]) begin out_Exp = in_Exp + 8'd48; out_Mant = in_Mant >> 48; end
        else if (in_Mant[174]) begin out_Exp = in_Exp + 8'd47; out_Mant = in_Mant >> 47; end
        else if (in_Mant[173]) begin out_Exp = in_Exp + 8'd46; out_Mant = in_Mant >> 46; end
        else if (in_Mant[172]) begin out_Exp = in_Exp + 8'd45; out_Mant = in_Mant >> 45; end
        else if (in_Mant[171]) begin out_Exp = in_Exp + 8'd44; out_Mant = in_Mant >> 44; end
        else if (in_Mant[170]) begin out_Exp = in_Exp + 8'd43; out_Mant = in_Mant >> 43; end
        else if (in_Mant[169]) begin out_Exp = in_Exp + 8'd42; out_Mant = in_Mant >> 42; end
        else if (in_Mant[168]) begin out_Exp = in_Exp + 8'd41; out_Mant = in_Mant >> 41; end
        else if (in_Mant[167]) begin out_Exp = in_Exp + 8'd40; out_Mant = in_Mant >> 40; end
        else if (in_Mant[166]) begin out_Exp = in_Exp + 8'd39; out_Mant = in_Mant >> 39; end
        else if (in_Mant[165]) begin out_Exp = in_Exp + 8'd38; out_Mant = in_Mant >> 38; end
        else if (in_Mant[164]) begin out_Exp = in_Exp + 8'd37; out_Mant = in_Mant >> 37; end
        else if (in_Mant[163]) begin out_Exp = in_Exp + 8'd36; out_Mant = in_Mant >> 36; end
        else if (in_Mant[162]) begin out_Exp = in_Exp + 8'd35; out_Mant = in_Mant >> 35; end
        else if (in_Mant[161]) begin out_Exp = in_Exp + 8'd34; out_Mant = in_Mant >> 34; end
        else if (in_Mant[160]) begin out_Exp = in_Exp + 8'd33; out_Mant = in_Mant >> 33; end
        else if (in_Mant[159]) begin out_Exp = in_Exp + 8'd32; out_Mant = in_Mant >> 32; end
        else if (in_Mant[158]) begin out_Exp = in_Exp + 8'd31; out_Mant = in_Mant >> 31; end
        else if (in_Mant[157]) begin out_Exp = in_Exp + 8'd30; out_Mant = in_Mant >> 30; end
        else if (in_Mant[156]) begin out_Exp = in_Exp + 8'd29; out_Mant = in_Mant >> 29; end
        else if (in_Mant[155]) begin out_Exp = in_Exp + 8'd28; out_Mant = in_Mant >> 28; end
        else if (in_Mant[154]) begin out_Exp = in_Exp + 8'd27; out_Mant = in_Mant >> 27; end
        else if (in_Mant[153]) begin out_Exp = in_Exp + 8'd26; out_Mant = in_Mant >> 26; end
        else if (in_Mant[152]) begin out_Exp = in_Exp + 8'd25; out_Mant = in_Mant >> 25; end
        else if (in_Mant[151]) begin out_Exp = in_Exp + 8'd24; out_Mant = in_Mant >> 24; end
        else if (in_Mant[150]) begin out_Exp = in_Exp + 8'd23; out_Mant = in_Mant >> 23; end
        else if (in_Mant[149]) begin out_Exp = in_Exp + 8'd22; out_Mant = in_Mant >> 22; end
        else if (in_Mant[148]) begin out_Exp = in_Exp + 8'd21; out_Mant = in_Mant >> 21; end
        else if (in_Mant[147]) begin out_Exp = in_Exp + 8'd20; out_Mant = in_Mant >> 20; end
        else if (in_Mant[146]) begin out_Exp = in_Exp + 8'd19; out_Mant = in_Mant >> 19; end
        else if (in_Mant[145]) begin out_Exp = in_Exp + 8'd18; out_Mant = in_Mant >> 18; end
        else if (in_Mant[144]) begin out_Exp = in_Exp + 8'd17; out_Mant = in_Mant >> 17; end
        else if (in_Mant[143]) begin out_Exp = in_Exp + 8'd16; out_Mant = in_Mant >> 16; end
        else if (in_Mant[142]) begin out_Exp = in_Exp + 8'd15; out_Mant = in_Mant >> 15; end
        else if (in_Mant[141]) begin out_Exp = in_Exp + 8'd14; out_Mant = in_Mant >> 14; end
        else if (in_Mant[140]) begin out_Exp = in_Exp + 8'd13; out_Mant = in_Mant >> 13; end
        else if (in_Mant[139]) begin out_Exp = in_Exp + 8'd12; out_Mant = in_Mant >> 12; end
        else if (in_Mant[138]) begin out_Exp = in_Exp + 8'd11; out_Mant = in_Mant >> 11; end
        else if (in_Mant[137]) begin out_Exp = in_Exp + 8'd10; out_Mant = in_Mant >> 10; end
        else if (in_Mant[136]) begin out_Exp = in_Exp + 8'd9; out_Mant = in_Mant >> 9; end
        else if (in_Mant[135]) begin out_Exp = in_Exp + 8'd8; out_Mant = in_Mant >> 8; end
        else if (in_Mant[134]) begin out_Exp = in_Exp + 8'd7; out_Mant = in_Mant >> 7; end
        else if (in_Mant[133]) begin out_Exp = in_Exp + 8'd6; out_Mant = in_Mant >> 6; end
        else if (in_Mant[132]) begin out_Exp = in_Exp + 8'd5; out_Mant = in_Mant >> 5; end
        else if (in_Mant[131]) begin out_Exp = in_Exp + 8'd4; out_Mant = in_Mant >> 4; end
        else if (in_Mant[130]) begin out_Exp = in_Exp + 8'd3; out_Mant = in_Mant >> 3; end
        else if (in_Mant[129]) begin out_Exp = in_Exp + 8'd2; out_Mant = in_Mant >> 2; end
        else if (in_Mant[128]) begin out_Exp = in_Exp + 8'd1; out_Mant = in_Mant >> 1; end
        else if (in_Mant[127]) begin out_Exp = in_Exp; out_Mant = in_Mant; end
        else if (in_Mant[126]) begin out_Exp = in_Exp - 8'd1; out_Mant = in_Mant << 1; end
        else if (in_Mant[125]) begin out_Exp = in_Exp - 8'd2; out_Mant = in_Mant << 2; end
        else if (in_Mant[124]) begin out_Exp = in_Exp - 8'd3; out_Mant = in_Mant << 3; end
        else if (in_Mant[123]) begin out_Exp = in_Exp - 8'd4; out_Mant = in_Mant << 4; end
        else if (in_Mant[122]) begin out_Exp = in_Exp - 8'd5; out_Mant = in_Mant << 5; end
        else if (in_Mant[121]) begin out_Exp = in_Exp - 8'd6; out_Mant = in_Mant << 6; end
        else if (in_Mant[120]) begin out_Exp = in_Exp - 8'd7; out_Mant = in_Mant << 7; end
        else if (in_Mant[119]) begin out_Exp = in_Exp - 8'd8; out_Mant = in_Mant << 8; end
        else if (in_Mant[118]) begin out_Exp = in_Exp - 8'd9; out_Mant = in_Mant << 9; end
        else if (in_Mant[117]) begin out_Exp = in_Exp - 8'd10; out_Mant = in_Mant << 10; end
        else if (in_Mant[116]) begin out_Exp = in_Exp - 8'd11; out_Mant = in_Mant << 11; end
        else if (in_Mant[115]) begin out_Exp = in_Exp - 8'd12; out_Mant = in_Mant << 12; end
        else if (in_Mant[114]) begin out_Exp = in_Exp - 8'd13; out_Mant = in_Mant << 13; end
        else if (in_Mant[113]) begin out_Exp = in_Exp - 8'd14; out_Mant = in_Mant << 14; end
        else if (in_Mant[112]) begin out_Exp = in_Exp - 8'd15; out_Mant = in_Mant << 15; end
        else if (in_Mant[111]) begin out_Exp = in_Exp - 8'd16; out_Mant = in_Mant << 16; end
        else if (in_Mant[110]) begin out_Exp = in_Exp - 8'd17; out_Mant = in_Mant << 17; end
        else if (in_Mant[109]) begin out_Exp = in_Exp - 8'd18; out_Mant = in_Mant << 18; end
        else if (in_Mant[108]) begin out_Exp = in_Exp - 8'd19; out_Mant = in_Mant << 19; end
        else if (in_Mant[107]) begin out_Exp = in_Exp - 8'd20; out_Mant = in_Mant << 20; end
        else if (in_Mant[106]) begin out_Exp = in_Exp - 8'd21; out_Mant = in_Mant << 21; end
        else if (in_Mant[105]) begin out_Exp = in_Exp - 8'd22; out_Mant = in_Mant << 22; end
        else if (in_Mant[104]) begin out_Exp = in_Exp - 8'd23; out_Mant = in_Mant << 23; end
        else if (in_Mant[103]) begin out_Exp = in_Exp - 8'd24; out_Mant = in_Mant << 24; end
        else if (in_Mant[102]) begin out_Exp = in_Exp - 8'd25; out_Mant = in_Mant << 25; end
        else if (in_Mant[101]) begin out_Exp = in_Exp - 8'd26; out_Mant = in_Mant << 26; end
        else if (in_Mant[100]) begin out_Exp = in_Exp - 8'd27; out_Mant = in_Mant << 27; end
        else if (in_Mant[99]) begin out_Exp = in_Exp - 8'd28; out_Mant = in_Mant << 28; end
        else if (in_Mant[98]) begin out_Exp = in_Exp - 8'd29; out_Mant = in_Mant << 29; end
        else if (in_Mant[97]) begin out_Exp = in_Exp - 8'd30; out_Mant = in_Mant << 30; end
        else if (in_Mant[96]) begin out_Exp = in_Exp - 8'd31; out_Mant = in_Mant << 31; end
        else if (in_Mant[95]) begin out_Exp = in_Exp - 8'd32; out_Mant = in_Mant << 32; end
        else if (in_Mant[94]) begin out_Exp = in_Exp - 8'd33; out_Mant = in_Mant << 33; end
        else if (in_Mant[93]) begin out_Exp = in_Exp - 8'd34; out_Mant = in_Mant << 34; end
        else if (in_Mant[92]) begin out_Exp = in_Exp - 8'd35; out_Mant = in_Mant << 35; end
        else if (in_Mant[91]) begin out_Exp = in_Exp - 8'd36; out_Mant = in_Mant << 36; end
        else if (in_Mant[90]) begin out_Exp = in_Exp - 8'd37; out_Mant = in_Mant << 37; end
        else if (in_Mant[89]) begin out_Exp = in_Exp - 8'd38; out_Mant = in_Mant << 38; end
        else if (in_Mant[88]) begin out_Exp = in_Exp - 8'd39; out_Mant = in_Mant << 39; end
        else if (in_Mant[87]) begin out_Exp = in_Exp - 8'd40; out_Mant = in_Mant << 40; end
        else if (in_Mant[86]) begin out_Exp = in_Exp - 8'd41; out_Mant = in_Mant << 41; end
        else if (in_Mant[85]) begin out_Exp = in_Exp - 8'd42; out_Mant = in_Mant << 42; end
        else if (in_Mant[84]) begin out_Exp = in_Exp - 8'd43; out_Mant = in_Mant << 43; end
        else if (in_Mant[83]) begin out_Exp = in_Exp - 8'd44; out_Mant = in_Mant << 44; end
        else if (in_Mant[82]) begin out_Exp = in_Exp - 8'd45; out_Mant = in_Mant << 45; end
        else if (in_Mant[81]) begin out_Exp = in_Exp - 8'd46; out_Mant = in_Mant << 46; end
        else if (in_Mant[80]) begin out_Exp = in_Exp - 8'd47; out_Mant = in_Mant << 47; end
        else if (in_Mant[79]) begin out_Exp = in_Exp - 8'd48; out_Mant = in_Mant << 48; end
        else if (in_Mant[78]) begin out_Exp = in_Exp - 8'd49; out_Mant = in_Mant << 49; end
        else if (in_Mant[77]) begin out_Exp = in_Exp - 8'd50; out_Mant = in_Mant << 50; end
        else if (in_Mant[76]) begin out_Exp = in_Exp - 8'd51; out_Mant = in_Mant << 51; end
        else if (in_Mant[75]) begin out_Exp = in_Exp - 8'd52; out_Mant = in_Mant << 52; end
        else if (in_Mant[74]) begin out_Exp = in_Exp - 8'd53; out_Mant = in_Mant << 53; end
        else if (in_Mant[73]) begin out_Exp = in_Exp - 8'd54; out_Mant = in_Mant << 54; end
        else if (in_Mant[72]) begin out_Exp = in_Exp - 8'd55; out_Mant = in_Mant << 55; end
        else if (in_Mant[71]) begin out_Exp = in_Exp - 8'd56; out_Mant = in_Mant << 56; end
        else if (in_Mant[70]) begin out_Exp = in_Exp - 8'd57; out_Mant = in_Mant << 57; end
        else if (in_Mant[69]) begin out_Exp = in_Exp - 8'd58; out_Mant = in_Mant << 58; end
        else if (in_Mant[68]) begin out_Exp = in_Exp - 8'd59; out_Mant = in_Mant << 59; end
        else if (in_Mant[67]) begin out_Exp = in_Exp - 8'd60; out_Mant = in_Mant << 60; end
        else if (in_Mant[66]) begin out_Exp = in_Exp - 8'd61; out_Mant = in_Mant << 61; end
        else if (in_Mant[65]) begin out_Exp = in_Exp - 8'd62; out_Mant = in_Mant << 62; end
        else if (in_Mant[64]) begin out_Exp = in_Exp - 8'd63; out_Mant = in_Mant << 63; end
        else if (in_Mant[63]) begin out_Exp = in_Exp - 8'd64; out_Mant = in_Mant << 64; end
        else if (in_Mant[62]) begin out_Exp = in_Exp - 8'd65; out_Mant = in_Mant << 65; end
        else if (in_Mant[61]) begin out_Exp = in_Exp - 8'd66; out_Mant = in_Mant << 66; end
        else if (in_Mant[60]) begin out_Exp = in_Exp - 8'd67; out_Mant = in_Mant << 67; end
        else if (in_Mant[59]) begin out_Exp = in_Exp - 8'd68; out_Mant = in_Mant << 68; end
        else if (in_Mant[58]) begin out_Exp = in_Exp - 8'd69; out_Mant = in_Mant << 69; end
        else if (in_Mant[57]) begin out_Exp = in_Exp - 8'd70; out_Mant = in_Mant << 70; end
        else if (in_Mant[56]) begin out_Exp = in_Exp - 8'd71; out_Mant = in_Mant << 71; end
        else if (in_Mant[55]) begin out_Exp = in_Exp - 8'd72; out_Mant = in_Mant << 72; end
        else if (in_Mant[54]) begin out_Exp = in_Exp - 8'd73; out_Mant = in_Mant << 73; end
        else if (in_Mant[53]) begin out_Exp = in_Exp - 8'd74; out_Mant = in_Mant << 74; end
        else if (in_Mant[52]) begin out_Exp = in_Exp - 8'd75; out_Mant = in_Mant << 75; end
        else if (in_Mant[51]) begin out_Exp = in_Exp - 8'd76; out_Mant = in_Mant << 76; end
        else if (in_Mant[50]) begin out_Exp = in_Exp - 8'd77; out_Mant = in_Mant << 77; end
        else if (in_Mant[49]) begin out_Exp = in_Exp - 8'd78; out_Mant = in_Mant << 78; end
        else if (in_Mant[48]) begin out_Exp = in_Exp - 8'd79; out_Mant = in_Mant << 79; end
        else if (in_Mant[47]) begin out_Exp = in_Exp - 8'd80; out_Mant = in_Mant << 80; end
        else if (in_Mant[46]) begin out_Exp = in_Exp - 8'd81; out_Mant = in_Mant << 81; end
        else if (in_Mant[45]) begin out_Exp = in_Exp - 8'd82; out_Mant = in_Mant << 82; end
        else if (in_Mant[44]) begin out_Exp = in_Exp - 8'd83; out_Mant = in_Mant << 83; end
        else if (in_Mant[43]) begin out_Exp = in_Exp - 8'd84; out_Mant = in_Mant << 84; end
        else if (in_Mant[42]) begin out_Exp = in_Exp - 8'd85; out_Mant = in_Mant << 85; end
        else if (in_Mant[41]) begin out_Exp = in_Exp - 8'd86; out_Mant = in_Mant << 86; end
        else if (in_Mant[40]) begin out_Exp = in_Exp - 8'd87; out_Mant = in_Mant << 87; end
        else if (in_Mant[39]) begin out_Exp = in_Exp - 8'd88; out_Mant = in_Mant << 88; end
        else if (in_Mant[38]) begin out_Exp = in_Exp - 8'd89; out_Mant = in_Mant << 89; end
        else if (in_Mant[37]) begin out_Exp = in_Exp - 8'd90; out_Mant = in_Mant << 90; end
        else if (in_Mant[36]) begin out_Exp = in_Exp - 8'd91; out_Mant = in_Mant << 91; end
        else if (in_Mant[35]) begin out_Exp = in_Exp - 8'd92; out_Mant = in_Mant << 92; end
        else if (in_Mant[34]) begin out_Exp = in_Exp - 8'd93; out_Mant = in_Mant << 93; end
        else if (in_Mant[33]) begin out_Exp = in_Exp - 8'd94; out_Mant = in_Mant << 94; end
        else if (in_Mant[32]) begin out_Exp = in_Exp - 8'd95; out_Mant = in_Mant << 95; end
        else if (in_Mant[31]) begin out_Exp = in_Exp - 8'd96; out_Mant = in_Mant << 96; end
        else if (in_Mant[30]) begin out_Exp = in_Exp - 8'd97; out_Mant = in_Mant << 97; end
        else if (in_Mant[29]) begin out_Exp = in_Exp - 8'd98; out_Mant = in_Mant << 98; end
        else if (in_Mant[28]) begin out_Exp = in_Exp - 8'd99; out_Mant = in_Mant << 99; end
        else if (in_Mant[27]) begin out_Exp = in_Exp - 8'd100; out_Mant = in_Mant << 100; end
        else if (in_Mant[26]) begin out_Exp = in_Exp - 8'd101; out_Mant = in_Mant << 101; end
        else if (in_Mant[25]) begin out_Exp = in_Exp - 8'd102; out_Mant = in_Mant << 102; end
        else if (in_Mant[24]) begin out_Exp = in_Exp - 8'd103; out_Mant = in_Mant << 103; end
        else if (in_Mant[23]) begin out_Exp = in_Exp - 8'd104; out_Mant = in_Mant << 104; end
        else if (in_Mant[22]) begin out_Exp = in_Exp - 8'd105; out_Mant = in_Mant << 105; end
        else if (in_Mant[21]) begin out_Exp = in_Exp - 8'd106; out_Mant = in_Mant << 106; end
        else if (in_Mant[20]) begin out_Exp = in_Exp - 8'd107; out_Mant = in_Mant << 107; end
        else if (in_Mant[19]) begin out_Exp = in_Exp - 8'd108; out_Mant = in_Mant << 108; end
        else if (in_Mant[18]) begin out_Exp = in_Exp - 8'd109; out_Mant = in_Mant << 109; end
        else if (in_Mant[17]) begin out_Exp = in_Exp - 8'd110; out_Mant = in_Mant << 110; end
        else if (in_Mant[16]) begin out_Exp = in_Exp - 8'd111; out_Mant = in_Mant << 111; end
        else if (in_Mant[15]) begin out_Exp = in_Exp - 8'd112; out_Mant = in_Mant << 112; end
        else if (in_Mant[14]) begin out_Exp = in_Exp - 8'd113; out_Mant = in_Mant << 113; end
        else if (in_Mant[13]) begin out_Exp = in_Exp - 8'd114; out_Mant = in_Mant << 114; end
        else if (in_Mant[12]) begin out_Exp = in_Exp - 8'd115; out_Mant = in_Mant << 115; end
        else if (in_Mant[11]) begin out_Exp = in_Exp - 8'd116; out_Mant = in_Mant << 116; end
        else if (in_Mant[10]) begin out_Exp = in_Exp - 8'd117; out_Mant = in_Mant << 117; end
        else if (in_Mant[9]) begin out_Exp = in_Exp - 8'd118; out_Mant = in_Mant << 118; end
        else if (in_Mant[8]) begin out_Exp = in_Exp - 8'd119; out_Mant = in_Mant << 119; end
        else if (in_Mant[7]) begin out_Exp = in_Exp - 8'd120; out_Mant = in_Mant << 120; end
        else if (in_Mant[6]) begin out_Exp = in_Exp - 8'd121; out_Mant = in_Mant << 121; end
        else if (in_Mant[5]) begin out_Exp = in_Exp - 8'd122; out_Mant = in_Mant << 122; end
        else if (in_Mant[4]) begin out_Exp = in_Exp - 8'd123; out_Mant = in_Mant << 123; end
        else if (in_Mant[3]) begin out_Exp = in_Exp - 8'd124; out_Mant = in_Mant << 124; end
        else if (in_Mant[2]) begin out_Exp = in_Exp - 8'd125; out_Mant = in_Mant << 125; end
        else if (in_Mant[1]) begin out_Exp = in_Exp - 8'd126; out_Mant = in_Mant << 126; end
        else begin out_Exp = in_Exp - 8'd127; out_Mant = in_Mant << 127; end
    end
endmodule