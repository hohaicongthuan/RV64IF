module Mant_Sqrt_Div_Ctrl(in_Clk, in_Rst_N, in_start, out_stall, out_load, out_shift_en);
    input   in_Clk, in_start, in_Rst_N;
    output  out_load, out_shift_en, out_stall;

    reg     [7:0] State_Reg;    // State register

    // Next-state Logics
    always @ (posedge in_Clk or negedge in_Rst_N) begin
        if (!in_Rst_N) begin
            State_Reg <= 0;
        end else begin
            case (State_Reg)
                8'd0: State_Reg <= (in_start) ? 8'd1 : 8'd0;
                8'd1: State_Reg <= 8'd2;
                8'd2: State_Reg <= 8'd3;
                8'd3: State_Reg <= 8'd4;
                8'd4: State_Reg <= 8'd5;
                8'd5: State_Reg <= 8'd6;
                8'd6: State_Reg <= 8'd7;
                8'd7: State_Reg <= 8'd8;
                8'd8: State_Reg <= 8'd9;
                8'd9: State_Reg <= 8'd10;
                8'd10: State_Reg <= 8'd11;
                8'd11: State_Reg <= 8'd12;
                8'd12: State_Reg <= 8'd13;
                8'd13: State_Reg <= 8'd14;
                8'd14: State_Reg <= 8'd15;
                8'd15: State_Reg <= 8'd16;
                8'd16: State_Reg <= 8'd17;
                8'd17: State_Reg <= 8'd18;
                8'd18: State_Reg <= 8'd19;
                8'd19: State_Reg <= 8'd20;
                8'd20: State_Reg <= 8'd21;
                8'd21: State_Reg <= 8'd22;
                8'd22: State_Reg <= 8'd23;
                8'd23: State_Reg <= 8'd24;
                8'd24: State_Reg <= 8'd25;
                8'd25: State_Reg <= 8'd26;
                8'd26: State_Reg <= 8'd27;
                8'd27: State_Reg <= 8'd28;
                8'd28: State_Reg <= 8'd29;
                8'd29: State_Reg <= 8'd30;
                8'd30: State_Reg <= 8'd31;
                8'd31: State_Reg <= 8'd32;
                8'd32: State_Reg <= 8'd33;
                8'd33: State_Reg <= 8'd34;
                8'd34: State_Reg <= 8'd35;
                8'd35: State_Reg <= 8'd36;
                8'd36: State_Reg <= 8'd37;
                8'd37: State_Reg <= 8'd38;
                8'd38: State_Reg <= 8'd39;
                8'd39: State_Reg <= 8'd40;
                8'd40: State_Reg <= 8'd41;
                8'd41: State_Reg <= 8'd42;
                8'd42: State_Reg <= 8'd43;
                8'd43: State_Reg <= 8'd44;
                8'd44: State_Reg <= 8'd45;
                8'd45: State_Reg <= 8'd46;
                8'd46: State_Reg <= 8'd47;
                8'd47: State_Reg <= 8'd48;
                8'd48: State_Reg <= 8'd49;
                8'd49: State_Reg <= 8'd50;
                8'd50: State_Reg <= 8'd51;
                8'd51: State_Reg <= 8'd52;
                8'd52: State_Reg <= 8'd53;
                8'd53: State_Reg <= 8'd54;
                8'd54: State_Reg <= 8'd55;
                8'd55: State_Reg <= 8'd56;
                8'd56: State_Reg <= 8'd57;
                8'd57: State_Reg <= 8'd58;
                8'd58: State_Reg <= 8'd59;
                8'd59: State_Reg <= 8'd60;
                8'd60: State_Reg <= 8'd61;
                8'd61: State_Reg <= 8'd62;
                8'd62: State_Reg <= 8'd63;
                8'd63: State_Reg <= 8'd64;
                8'd64: State_Reg <= 8'd65;
                8'd65: State_Reg <= 8'd66;
                8'd66: State_Reg <= 8'd67;
                8'd67: State_Reg <= 8'd68;
                8'd68: State_Reg <= 8'd69;
                8'd69: State_Reg <= 8'd70;
                8'd70: State_Reg <= 8'd71;
                8'd71: State_Reg <= 8'd72;
                8'd72: State_Reg <= 8'd73;
                8'd73: State_Reg <= 8'd74;
                8'd74: State_Reg <= 8'd75;
                8'd75: State_Reg <= 8'd76;
                8'd76: State_Reg <= 8'd77;
                8'd77: State_Reg <= 8'd78;
                8'd78: State_Reg <= 8'd79;
                8'd79: State_Reg <= 8'd80;
                8'd80: State_Reg <= 8'd81;
                8'd81: State_Reg <= 8'd82;
                8'd82: State_Reg <= 8'd83;
                8'd83: State_Reg <= 8'd84;
                8'd84: State_Reg <= 8'd85;
                8'd85: State_Reg <= 8'd86;
                8'd86: State_Reg <= 8'd87;
                8'd87: State_Reg <= 8'd88;
                8'd88: State_Reg <= 8'd89;
                8'd89: State_Reg <= 8'd90;
                8'd90: State_Reg <= 8'd91;
                8'd91: State_Reg <= 8'd92;
                8'd92: State_Reg <= 8'd93;
                8'd93: State_Reg <= 8'd94;
                8'd94: State_Reg <= 8'd95;
                8'd95: State_Reg <= 8'd96;
                8'd96: State_Reg <= 8'd97;
                8'd97: State_Reg <= 8'd98;
                8'd98: State_Reg <= 8'd99;
                8'd99: State_Reg <= 8'd100;
                8'd100: State_Reg <= 8'd101;
                8'd101: State_Reg <= 8'd102;
                8'd102: State_Reg <= 8'd103;
                8'd103: State_Reg <= 8'd104;
                8'd104: State_Reg <= 8'd105;
                8'd105: State_Reg <= 8'd106;
                8'd106: State_Reg <= 8'd107;
                8'd107: State_Reg <= 8'd108;
                8'd108: State_Reg <= 8'd109;
                8'd109: State_Reg <= 8'd110;
                8'd110: State_Reg <= 8'd111;
                8'd111: State_Reg <= 8'd112;
                8'd112: State_Reg <= 8'd113;
                8'd113: State_Reg <= 8'd114;
                8'd114: State_Reg <= 8'd115;
                8'd115: State_Reg <= 8'd116;
                8'd116: State_Reg <= 8'd117;
                8'd117: State_Reg <= 8'd118;
                8'd118: State_Reg <= 8'd119;
                8'd119: State_Reg <= 8'd120;
                8'd120: State_Reg <= 8'd121;
                8'd121: State_Reg <= 8'd122;
                8'd122: State_Reg <= 8'd123;
                8'd123: State_Reg <= 8'd124;
                8'd124: State_Reg <= 8'd125;
                8'd125: State_Reg <= 8'd126;
                8'd126: State_Reg <= 8'd127;
                8'd127: State_Reg <= 8'd128;
                8'd128: State_Reg <= 8'd129;
                8'd129: State_Reg <= 8'd130;
                8'd130: State_Reg <= 8'd131;
                8'd131: State_Reg <= 8'd132;
                8'd132: State_Reg <= 8'd133;
                8'd133: State_Reg <= 8'd134;
                8'd134: State_Reg <= 8'd135;
                8'd135: State_Reg <= 8'd136;
                8'd136: State_Reg <= 8'd137;
                8'd137: State_Reg <= 8'd138;
                8'd138: State_Reg <= 8'd139;
                8'd139: State_Reg <= 8'd140;
                8'd140: State_Reg <= 8'd141;
                8'd141: State_Reg <= 8'd142;
                8'd142: State_Reg <= 8'd143;
                8'd143: State_Reg <= 8'd144;
                8'd144: State_Reg <= 8'd145;
                8'd145: State_Reg <= 8'd146;
                8'd146: State_Reg <= 8'd147;
                8'd147: State_Reg <= 8'd148;
                8'd148: State_Reg <= 8'd149;
                8'd149: State_Reg <= 8'd150;
                8'd150: State_Reg <= 8'd151;
                8'd151: State_Reg <= 8'd152;
                8'd152: State_Reg <= 8'd153;
                8'd153: State_Reg <= 8'd154;
                8'd154: State_Reg <= 8'd155;
                8'd155: State_Reg <= 8'd156;
                8'd156: State_Reg <= 8'd157;
                8'd157: State_Reg <= 8'd158;
                8'd158: State_Reg <= 8'd159;
                8'd159: State_Reg <= 8'd160;
                8'd160: State_Reg <= 8'd161;
                8'd161: State_Reg <= 8'd162;
                8'd162: State_Reg <= 8'd163;
                8'd163: State_Reg <= 8'd164;
                8'd164: State_Reg <= 8'd165;
                8'd165: State_Reg <= 8'd166;
                8'd166: State_Reg <= 8'd167;
                8'd167: State_Reg <= 8'd168;
                8'd168: State_Reg <= 8'd169;
                8'd169: State_Reg <= 8'd170;
                8'd170: State_Reg <= 8'd171;
                8'd171: State_Reg <= 8'd172;
                8'd172: State_Reg <= 8'd173;
                8'd173: State_Reg <= 8'd174;
                8'd174: State_Reg <= 8'd175;
                8'd175: State_Reg <= 8'd176;
                8'd176: State_Reg <= 8'd177;
                8'd177: State_Reg <= 8'd178;
                8'd178: State_Reg <= 8'd179;
                8'd179: State_Reg <= 8'd180;
                8'd180: State_Reg <= 8'd181;
                8'd181: State_Reg <= 8'd182;
                8'd182: State_Reg <= 8'd183;
                8'd183: State_Reg <= 8'd184;
                8'd184: State_Reg <= 8'd185;
                8'd185: State_Reg <= 8'd186;
                8'd186: State_Reg <= 8'd187;
                8'd187: State_Reg <= 8'd188;
                8'd188: State_Reg <= 8'd189;
                8'd189: State_Reg <= 8'd190;
                8'd190: State_Reg <= 8'd191;
                8'd191: State_Reg <= 8'd192;
                8'd192: State_Reg <= 8'd193;
                8'd193: State_Reg <= 8'd194;
                8'd194: State_Reg <= 8'd195;
                8'd195: State_Reg <= 8'd196;
                8'd196: State_Reg <= 8'd197;
                8'd197: State_Reg <= 8'd198;
                8'd198: State_Reg <= 8'd199;
                8'd199: State_Reg <= 8'd200;
                8'd200: State_Reg <= 8'd201;
                8'd201: State_Reg <= 8'd202;
                8'd202: State_Reg <= 8'd203;
                8'd203: State_Reg <= 8'd204;
                8'd204: State_Reg <= 8'd205;
                8'd205: State_Reg <= 8'd206;
                8'd206: State_Reg <= 8'd207;
                8'd207: State_Reg <= 8'd208;
                8'd208: State_Reg <= 8'd209;
                8'd209: State_Reg <= 8'd210;
                8'd210: State_Reg <= 8'd211;
                8'd211: State_Reg <= 8'd212;
                8'd212: State_Reg <= 8'd213;
                8'd213: State_Reg <= 8'd214;
                8'd214: State_Reg <= 8'd215;
                8'd215: State_Reg <= 8'd216;
                8'd216: State_Reg <= 8'd217;
                8'd217: State_Reg <= 8'd218;
                8'd218: State_Reg <= 8'd219;
                8'd219: State_Reg <= 8'd220;
                8'd220: State_Reg <= 8'd221;
                8'd221: State_Reg <= 8'd222;
                8'd222: State_Reg <= 8'd223;
                8'd223: State_Reg <= 8'd224;
                8'd224: State_Reg <= 8'd225;
                8'd225: State_Reg <= 8'd226;
                8'd226: State_Reg <= 8'd227;
                8'd227: State_Reg <= 8'd228;
                8'd228: State_Reg <= 8'd229;
                8'd229: State_Reg <= 8'd230;
                8'd230: State_Reg <= 8'd231;
                8'd231: State_Reg <= 8'd232;
                8'd232: State_Reg <= 8'd233;
                8'd233: State_Reg <= 8'd234;
                8'd234: State_Reg <= 8'd235;
                8'd235: State_Reg <= 8'd236;
                8'd236: State_Reg <= 8'd237;
                8'd237: State_Reg <= 8'd238;
                8'd238: State_Reg <= 8'd239;
                8'd239: State_Reg <= 8'd240;
                8'd240: State_Reg <= 8'd241;
                8'd241: State_Reg <= 8'd242;
                8'd242: State_Reg <= 8'd243;
                8'd243: State_Reg <= 8'd244;
                8'd244: State_Reg <= 8'd245;
                8'd245: State_Reg <= 8'd246;
                8'd246: State_Reg <= 8'd247;
                8'd247: State_Reg <= 8'd248;
                8'd248: State_Reg <= 8'd249;
                8'd249: State_Reg <= 8'd250;
                8'd250: State_Reg <= 8'd251;
                8'd251: State_Reg <= 8'd252;
                8'd252: State_Reg <= 8'd253;
                8'd253: State_Reg <= 8'd254;
                8'd254: State_Reg <= 8'd255;
                8'd255: State_Reg <= 8'd0;
                default: State_Reg <= 8'd0;
            endcase
        end
    end

    // Output logics
    assign out_load     = (State_Reg == 8'd1) ? 1'b1 : 1'b0;
    assign out_shift_en = (State_Reg == 8'd0 | State_Reg == 8'd255) ? 1'b0 : 1'b1;
    assign out_stall    = (State_Reg < 8'd255 & in_start) ? 1'b1 : 1'b0;
endmodule